/*
 *  picoSoC_hardware -- SoC Hardware for RISCV-32I core.
 *
 *  Copyright (C) 2021-2021 Junnan Li <lijunnan@nudt.edu.cn>.
 *  Copyright and related rights are licensed under the MIT license.
 *
 *  Data: 2021.12.03
 *  Description: This module is used to connect Pico_top and configuration.
 */

module um_for_cpu(
  input               clk,
  input               rst_n,
    
  input               data_in_valid,
  input       [133:0] data_in,  // 2'b01 is head, 2'b00 is body, and 2'b10 is tail;
  
  output reg          data_out_valid,
  output reg  [133:0] data_out,

  //* left for packet process;
  output wire         mem_wren,
  output wire         mem_rden,
  output wire [31:0]  mem_addr,
  output wire [31:0]  mem_wdata,
  input       [31:0]  mem_rdata,
  output wire         cpu_ready
);

  /** TODO:*/

  (* mark_debug = "true"*)wire          conf_rden, conf_wren;
  (* mark_debug = "true"*)wire [31:0]   conf_addr, conf_wdata, conf_rdata;
  (* mark_debug = "true"*)wire          conf_sel;
  (* mark_debug = "true"*)wire          print_valid;
  (* mark_debug = "true"*)wire [7:0]    print_value;
  (* mark_debug = "true"*)wire          data_valid_confMem;
  (* mark_debug = "true"*)wire [133:0]  data_confMem;
  // fifo interface
  reg           rdreq_pkt;
  wire [133:0]  q_pkt;
  reg  [7:0]    count_pkt;  // number of packet in the fifo;
  
  assign cpu_ready  = 1'b1;
  assign mem_wren   = 1'b0;
  assign mem_rden   = 1'b0;
  assign mem_addr   = 32'b0;
  assign mem_wdata  = 32'b0;

  Pico_top picoTop(
    .clk(clk),
    .resetn(rst_n),

    .conf_rden(conf_rden),
    .conf_wren(conf_wren),
    .conf_addr(conf_addr),
    .conf_wdata(conf_wdata),
    .conf_rdata(conf_rdata),
    .conf_sel(conf_sel),

    .print_valid(print_valid),
    .print_value(print_value)
  );

  conf_mem confMem(
    .clk(clk),
    .resetn(rst_n),

    .data_in_valid(data_in_valid),
    .data_in(data_in),
    .data_out_valid(data_valid_confMem),
    .data_out(data_confMem),

    .conf_rden(conf_rden),
    .conf_wren(conf_wren),
    .conf_addr(conf_addr),
    .conf_wdata(conf_wdata),
    .conf_rdata(conf_rdata),
    .conf_sel(conf_sel),

    .print_valid(print_valid),
    .print_value(print_value)
  );


  /** fifo used to store packet generated by cpu*/
  fifo_134b_512 pkt_buffer(
    .clk(clk),
    .srst(!rst_n),
    .din(data_confMem),
    .wr_en(data_valid_confMem),
    .rd_en(rdreq_pkt),
    .dout(q_pkt),
    .full(),
    .empty()
  );

  /** output packet */
  reg         state_out;
  localparam  IDLE_S      = 1'b0,
              READ_FIFO_S = 1'b1;
  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      // reset
      count_pkt       <= 8'b0;
      // output packet;
      state_out       <= IDLE_S;
      data_out_valid  <= 1'b0;
      data_out        <= 134'b0;
      rdreq_pkt       <= 1'b0;
    end
    else begin
      //* count packets;
      if((data_confMem[133:132] == 2'b10 && data_valid_confMem == 1'b1) &&
        (data_out[133:132] == 2'b01 && data_out_valid == 1'b1))
          count_pkt   <= count_pkt;
      else if(data_confMem[133:132] == 2'b10 && data_valid_confMem == 1'b1)
        count_pkt     <= count_pkt + 8'd1;
      else if(data_out[133:132] == 2'b01 && data_out_valid == 1'b1)
        count_pkt     <= count_pkt - 8'd1;
      else
        count_pkt     <= count_pkt;

      (* full_case *)
      case(state_out)
        IDLE_S: begin
          data_out_valid  <= 1'b0;
          if(count_pkt != 0) begin
            rdreq_pkt     <= 1'b1;
            state_out     <= READ_FIFO_S;
          end
          else begin
            rdreq_pkt     <= 1'b0;
            state_out     <= IDLE_S;
          end
        end
        READ_FIFO_S: begin
          data_out_valid  <= 1'b1;
          data_out        <= q_pkt;
          if(q_pkt[133:132] == 2'b10) begin
            rdreq_pkt     <= 1'b0;
            state_out     <= IDLE_S;
          end
          else begin
            rdreq_pkt     <= 1'b1;
            state_out     <= READ_FIFO_S;
          end
        end
      endcase 
    end
  end

  
endmodule    
